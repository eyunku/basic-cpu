// Goku's D-flipflop

// simple dff
module dff (q, d, wen, clk, rst);
    output q; //DFF output
    input d; //DFF input
    input wen; //Write Enable
    input clk; //Clock
    input rst; //Reset (used synchronously)

    reg state;

    assign q = state;

    always @(posedge clk) begin
    state <= rst ? 0 : (wen ? d : state);
    end
endmodule
