module t_integration_Controller_Arbitration():
    
endmodule